module add_one()
