module mixer(CLOCK_50, 
						 audio0,
						 audio1,
						 audio2,
						 audio3,
						 audio4,
						 audio5,
						 audio6,
						 audio7);
	input CLOCK_50;
	input [15:0] ;


endmodule
