module triangle_wave #(parameter ACCUMULATOR_BITS = 24,
											 parameter OUTPUT_BITS = 12)
	(input [ACCUMULATOR_BITS-1:0] accumulator,
	 output wire [OUTPUT_BITS-1:0] out,
	 input en_ringmod,
	 input ringmod_source
	 );

	 

endmodule