module synth_snare();



endmodule
