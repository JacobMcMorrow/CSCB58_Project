module synth_snare();

	// Oscilator section
	// Sine 180Hz

	// Sine 330Hz

	// Triangle 111Hz

	// Freq shift triangle 

	// 

	// Noise section
	//

	
	// Out mixer
	

endmodule
